/opt/cadence/FreePDK45/osu_soc/lib/files/gscl45nm.lef